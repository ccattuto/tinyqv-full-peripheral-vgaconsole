// Synthesis-friendly: explicit array init + indexed combinational read.
module char_rom #(
    parameter DATA_WIDTH = 35,     // 35 bits per character
    parameter ADDR_WIDTH = 7,      // address width
    parameter ADDR_MIN   = 32,
    parameter ADDR_MAX   = 127
)(
    input  wire [ADDR_WIDTH-1:0] address,
    output wire [DATA_WIDTH-1:0] data
);

reg [DATA_WIDTH-1:0] d;

// bit permutation (unchanged)
assign data = { d[32], d[24], d[21], d[26], d[19], d[29], d[17], d[13], d[25], d[12],
                d[0],  d[14], d[4],  d[28], d[18], d[3],  d[31], d[22], d[1],  d[11],
                d[34], d[15], d[30], d[23], d[2],  d[8],  d[27], d[7],  d[33], d[20],
                d[10], d[9],  d[5],  d[16], d[6] };

// ROM storage: addresses 32..127
reg [DATA_WIDTH-1:0] mem [ADDR_MIN:ADDR_MAX];

initial begin
    mem[7'd32]  = 35'b00000000000000000000000000000000000;
    mem[7'd33]  = 35'b00001000000011000000000000010110000;
    mem[7'd34]  = 35'b01000001000100000011000001000000000;
    mem[7'd35]  = 35'b11011011111100001111100001000010111;
    mem[7'd36]  = 35'b01011001010011000100011000110110111;
    mem[7'd37]  = 35'b01100110001010100111001000101000000;
    mem[7'd38]  = 35'b00101000100001101110001000010010111;
    mem[7'd39]  = 35'b00001001000000000000000001010100010;
    mem[7'd40]  = 35'b00000010001100000000010001010000010;
    mem[7'd41]  = 35'b00010000100000000011110000010000000;
    mem[7'd42]  = 35'b00011110000111100001111100110111010;
    mem[7'd43]  = 35'b00011000000010000000010100010011010;
    mem[7'd44]  = 35'b00000000000001000100110000000010000;
    mem[7'd45]  = 35'b00010000000010000000000100000001010;
    mem[7'd46]  = 35'b00000000001001000100010000000000000;
    mem[7'd47]  = 35'b00000010000010000001001000100000000;
    mem[7'd48]  = 35'b10000110101011101011001101100101101;
    mem[7'd49]  = 35'b01001000101011000000010000010110000;
    mem[7'd50]  = 35'b10110000101011111010001001100100010;
    mem[7'd51]  = 35'b00010100101011000011001011101100001;
    mem[7'd52]  = 35'b00010011001100001101100101010010001;
    mem[7'd53]  = 35'b00001100101101100011001011001101101;
    mem[7'd54]  = 35'b01010100101011001000001111000100111;
    mem[7'd55]  = 35'b10010000010000010010000011101110000;
    mem[7'd56]  = 35'b10010100101011101010001001100100111;
    mem[7'd57]  = 35'b10010000100011110110000001100101111;
    mem[7'd58]  = 35'b00001000000000000000000000000010000;
    mem[7'd59]  = 35'b00001000100000000000010000000010000;
    mem[7'd60]  = 35'b00101001000000000100000010000010010;
    mem[7'd61]  = 35'b10001010000100001001100000000010101;
    mem[7'd62]  = 35'b00000000100000000011110000010001000;
    mem[7'd63]  = 35'b10010000000011100010000001100110000;
    mem[7'd64]  = 35'b10111000101011101010101101100111100;
    mem[7'd65]  = 35'b11100111000000011000101100000111101;
    mem[7'd66]  = 35'b10010100101011111010001101101100111;
    mem[7'd67]  = 35'b00000100101001101010001101100100100;
    mem[7'd68]  = 35'b10000100101001111010001101101101101;
    mem[7'd69]  = 35'b00110000101011111010001111001100110;
    mem[7'd70]  = 35'b00010000000010111010001111001100110;
    mem[7'd71]  = 35'b00100100101001101010101111100100101;
    mem[7'd72]  = 35'b10110100000010111000001110101001111;
    mem[7'd73]  = 35'b00001000101011000010010001010110000;
    mem[7'd74]  = 35'b00010001100001000101101011000100000;
    mem[7'd75]  = 35'b00101001000000111100001110001010110;
    mem[7'd76]  = 35'b00100000101001111000001100001000100;
    mem[7'd77]  = 35'b11101101000010111000001110101011101;
    mem[7'd78]  = 35'b10100100000110111000101110101001101;
    mem[7'd79]  = 35'b10000100101001101010001101100101101;
    mem[7'd80]  = 35'b10010000000010111010001101101100110;
    mem[7'd81]  = 35'b10100000100001101110001101100111101;
    mem[7'd82]  = 35'b10110000000010111110001101101110110;
    mem[7'd83]  = 35'b00010100101011100010001001100100111;
    mem[7'd84]  = 35'b00001000000011100010010011111110000;
    mem[7'd85]  = 35'b10000100101001101000001110101001101;
    mem[7'd86]  = 35'b10000000010001101100000110101001101;
    mem[7'd87]  = 35'b10000100101010101000011110101011101;
    mem[7'd88]  = 35'b00100110000110110001101010101000000;
    mem[7'd89]  = 35'b00000000000111100001010010101010000;
    mem[7'd90]  = 35'b00110010101011010011001011101100010;
    mem[7'd91]  = 35'b01100010111101000010000011000100010;
    mem[7'd92]  = 35'b00000100000110100000100000000000000;
    mem[7'd93]  = 35'b10100100101001000010000011100101001;
    mem[7'd94]  = 35'b11000001000000000000000000000100100;
    mem[7'd95]  = 35'b00100000101001010000000000000000000;
    mem[7'd96]  = 35'b01011000000000000010000000010100000;
    mem[7'd97]  = 35'b00111010101101000100101000000010000;
    mem[7'd98]  = 35'b00001100011001111001001100001001111;
    mem[7'd99]  = 35'b00001100101101001001001100000001000;
    mem[7'd100] = 35'b10111100100101001100001110100001001;
    mem[7'd101] = 35'b00001010101101001001101100000011001;
    mem[7'd102] = 35'b00011000000011000000010001110010010;
    mem[7'd103] = 35'b00111100010100001001110100000001001;
    mem[7'd104] = 35'b00101100000000111001001100001001111;
    mem[7'd105] = 35'b00001000101111000000010000000110000;
    mem[7'd106] = 35'b00010000100001000101101001000000000;
    mem[7'd107] = 35'b00000010001010111001011100001000100;
    mem[7'd108] = 35'b00001000101011000010010000010110000;
    mem[7'd109] = 35'b00100100000111011001011100000011101;
    mem[7'd110] = 35'b00101100000000011001001100000001111;
    mem[7'd111] = 35'b00001100101101001001001100000001001;
    mem[7'd112] = 35'b00001010000000011101011100000001111;
    mem[7'd113] = 35'b10111100010100001000110100000001001;
    mem[7'd114] = 35'b00001000000000011001001100000001110;
    mem[7'd115] = 35'b10001110101101010001100100000010000;
    mem[7'd116] = 35'b10001100001110000001010000010110100;
    mem[7'd117] = 35'b10100100100001001100001100000001101;
    mem[7'd118] = 35'b10000000010001001100000100000001101;
    mem[7'd119] = 35'b10000100101000001000011100000011101;
    mem[7'd120] = 35'b10110000010000010100000000000010110;
    mem[7'd121] = 35'b10100110000000010000100100000011101;
    mem[7'd122] = 35'b10111000111101010001000000000010100;
    mem[7'd123] = 35'b00001000001000000000010001010010010;
    mem[7'd124] = 35'b00001000000001000000010000010110000;
    mem[7'd125] = 35'b00011000100000000010010000010010000;
    mem[7'd126] = 35'b00000000000000100011000000110000000;
    mem[7'd127] = 35'b11111111111111111111111111111111111;
end

// Combinational indexed read with range guard
always @* begin
  if (address >= ADDR_MIN)
    d = mem[address];
  else
    d = {DATA_WIDTH{1'b1}}; // default = all ones (Verilog-2001 portable)
end

endmodule
