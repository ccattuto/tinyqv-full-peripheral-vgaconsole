/*
 * Copyright (c) 2025 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

// Change the name of this module to something that reflects its functionality and includes your name for uniqueness
// For example tqvp_yourname_spi for an SPI peripheral.
// Then edit tt_wrapper.v line 41 and change tqvp_example to your chosen module name.
module tqvp_example (
    input         clk,          // Clock - the TinyQV project clock is normally set to 64MHz.
    input         rst_n,        // Reset_n - low to reset.

    input  [7:0]  ui_in,        // The input PMOD, always available.  Note that ui_in[7] is normally used for UART RX.
                                // The inputs are synchronized to the clock, note this will introduce 2 cycles of delay on the inputs.

    output [7:0]  uo_out,       // The output PMOD.  Each wire is only connected if this peripheral is selected.
                                // Note that uo_out[0] is normally used for UART TX.

    input [5:0]   address,      // Address within this peripheral's address space
    input [31:0]  data_in,      // Data in to the peripheral, bottom 8, 16 or all 32 bits are valid on write.

    // Data read and write requests from the TinyQV core.
    input [1:0]   data_write_n, // 11 = no write, 00 = 8-bits, 01 = 16-bits, 10 = 32-bits
    input [1:0]   data_read_n,  // 11 = no read,  00 = 8-bits, 01 = 16-bits, 10 = 32-bits
    
    output [31:0] data_out,     // Data out from the peripheral, bottom 8, 16 or all 32 bits are valid on read when data_ready is high.
    output        data_ready,

    output        user_interrupt  // Dedicated interrupt request for this peripheral
);

    localparam NUM_ROWS = 3;
    localparam NUM_COLS = 10;
    localparam NUM_CHARS = NUM_ROWS * NUM_COLS;
    localparam ROWS_ADDR_WIDTH = $clog2(NUM_ROWS);
    localparam COLS_ADDR_WIDTH = $clog2(NUM_COLS);
    localparam CHARS_ADDR_WIDTH = $clog2(NUM_CHARS);

    // Text buffer (7-bit chars)
    reg [6:0] text[0:NUM_CHARS-1];
    reg [5:0] text_color[0:NUM_CHARS-1];
    reg [5:0] bg_color;

    // ----- HOST INTERFACE -----
    
    // Writes to memory-mapped text buffer: only write lowest 8 bits
    always @(posedge clk) begin
        if (!rst_n) begin
            bg_color <= 6'b010000;
        end else begin
            if (address < NUM_CHARS) begin
                if (data_write_n != 2'b11) begin
                    text[address[CHARS_ADDR_WIDTH-1:0]] <= data_in[6:0];
                end
                if (data_write_n == 2'b00) begin
                    text_color[address[CHARS_ADDR_WIDTH-1:0]] <= 6'b011100;     // default text color
                end else if (data_write_n != 2'b11) begin
                    text_color[address[CHARS_ADDR_WIDTH-1:0]] <= data_in[13:8]; // set color
                end
            end else if (address == 6'h3F && data_write_n != 2'b11) begin
                bg_color <= data_in[5:0];
            end
        end
    end

    // Register reads
    assign data_out = (address < NUM_CHARS) ? {18'h0, text_color[address[CHARS_ADDR_WIDTH-1:0]], 1'b0, text[address[CHARS_ADDR_WIDTH-1:0]]} : (address == 6'h3F) ? {26'h0, bg_color} : 32'h0;

    // All reads complete in 1 clock
    assign data_ready = 1;

    // No interrupt handling
    assign user_interrupt = 0;

    wire _unused = &{data_read_n, 1'b0};


    // ----- VGA INTERFACE -----

    localparam VGA_WIDTH = 640;
    localparam VGA_HEIGHT = 480;
    localparam VGA_FRAME_XMIN = 80;
    localparam VGA_FRAME_XMAX = VGA_WIDTH - 80;
    localparam VGA_FRAME_YMIN = 128;
    localparam VGA_FRAME_YMAX = VGA_HEIGHT - 160;

    // VGA signals
    wire hsync;
    wire vsync;
    wire [1:0] R;
    wire [1:0] G;
    wire [1:0] B;
    wire video_active;
    wire [9:0] pix_x;
    wire [9:0] pix_y;

    // TinyVGA PMOD
    assign uo_out = {hsync, B[0], G[0], R[0], vsync, B[1], G[1], R[1]};

    hvsync_generator hvsync_gen(
        .clk(clk),
        .reset(~rst_n),
        .hsync(hsync),
        .vsync(vsync),
        .display_on(video_active),
        .hpos(pix_x),
        .vpos(pix_y)
    );

    wire frame_active;
    assign frame_active = (pix_x >= VGA_FRAME_XMIN && pix_x < VGA_FRAME_XMAX && pix_y >= VGA_FRAME_YMIN && pix_y < VGA_FRAME_YMAX) ? 1 : 0;

    // (x,y) coordinates relative to frame
    wire [9:0] pix_x_frame, pix_y_frame;
    assign pix_x_frame = pix_x - VGA_FRAME_XMIN;
    assign pix_y_frame = pix_y - VGA_FRAME_YMIN;

    // Character pixels are 8x8 squares in the VGA frame.
    // Character glyphs are 5x7 and padded in a 6x8 character box.

    // (x,y) character coordinates in NUM_ROWS x NUM_COLS text buffer
    wire [COLS_ADDR_WIDTH-1:0] char_x;
    wire [ROWS_ADDR_WIDTH-1:0] char_y;
    assign char_x = (pix_x_frame / 6) >> 3; // divide by 48 (VGA char width is 48 pixels)
    assign char_y = pix_y_frame >> 6;       // divide by 64 (VGA char height is 64 pixels)

    // Drive character ROM input
    wire [6:0] char_index;
    assign char_index = text[char_y * NUM_COLS + char_x];

    // Character color
    wire [5:0] char_color;
    assign char_color = text_color[char_y * NUM_COLS + char_x];

    // Character pixel coordinates relative to the 5x7 glyph padded in a 6x8 character box
    wire [2:0] rel_x;
    wire [2:0] rel_y;
    assign rel_x = pix_x_frame[9:3] % 6;    // remainder of division by 6
    assign rel_y = pix_y_frame[9:3] & 7;    // remainder of division by 8

    // Character pixel index in the 35-bit wide character ROM (rel_y * 5 + rel_x)
    wire [5:0] offset;
    assign offset = (rel_y << 2) + rel_y + rel_x;

    // Look up character pixel value in character ROM,
    // handling 1-pixel padding along x and y directions.
    wire char_pixel;
    assign char_pixel = ((rel_y == 7) || (rel_x == 5)) ? 0 : char_data[offset];

    // generate RGB signals
    wire pixel_on;
    assign pixel_on = frame_active & char_pixel;
    assign R = ~video_active ? 2'b00 : (pixel_on ? char_color[1:0] : bg_color[1:0]);
    assign G = ~video_active ? 2'b00 : (pixel_on ? char_color[3:2] : bg_color[3:2]);
    assign B = ~video_active ? 2'b00 : (pixel_on ? char_color[5:4] : bg_color[5:4]);

    // ----- CHARACTER ROM -----

    wire [34:0] char_data;

    char_rom char_rom_inst (
        .address(char_index),
        .data(char_data) 
    );

endmodule
